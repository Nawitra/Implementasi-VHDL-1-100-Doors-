LIBRARY IEEE  ; 
LIBRARY STD  ; 
USE IEEE.STD_LOGIC_1164.ALL  ; 
USE IEEE.STD_LOGIC_TEXTIO.ALL  ; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL  ; 
USE STD.TEXTIO.ALL  ; 
ENTITY TESTBENCH_PINTU  IS 
END ; 
 
ARCHITECTURE TESTBENCH_PINTU_ARCH OF TESTBENCH_PINTU IS
  SIGNAL OUTPUT   :  STD_LOGIC_VECTOR (1 TO 100) := (OTHERS =>  '0')  ; 
  SIGNAL RST   :  STD_LOGIC  ; 
  SIGNAL CLK   :  STD_LOGIC  ; 
  COMPONENT DOORS  
    PORT ( 
      OUTPUT  : INOUT STD_LOGIC_VECTOR (1 TO 100) ; 
      RST  : IN STD_LOGIC ; 
      CLK  : IN STD_LOGIC ); 
  END COMPONENT ; 
BEGIN
  DUT  : DOORS  
    PORT MAP ( 
      OUTPUT   => OUTPUT  ,
      RST   => RST  ,
      CLK   => CLK   ) ; 



-- "CLOCK PATTERN" : DUTYCYCLE = 50
-- START TIME = 0 PS, END TIME = 1 NS, PERIOD = 100 PS
  PROCESS
	BEGIN
	 CLK  <= '0'  ;
	WAIT FOR 50 PS ;
-- 50 PS, SINGLE LOOP TILL START PERIOD.
	FOR Z IN 1 TO 9
	LOOP
	    CLK  <= '1'  ;
	   WAIT FOR 50 PS ;
	    CLK  <= '0'  ;
	   WAIT FOR 50 PS ;
-- 950 PS, REPEAT PATTERN IN LOOP.
	END  LOOP;
	 CLK  <= '1'  ;
	WAIT FOR 50 PS ;
-- DUMPED VALUES TILL 1 NS
	WAIT;
 END PROCESS;


-- "CONSTANT PATTERN"
-- START TIME = 50 PS, END TIME = 10 NS, PERIOD = 0 PS
  PROCESS
	BEGIN
	 RST  <= '1'  ;
	WAIT FOR 50 PS ;
	 RST  <= '0'  ;
	WAIT FOR 9950 PS ;
-- DUMPED VALUES TILL 10 NS
	WAIT;
 END PROCESS;
END;
